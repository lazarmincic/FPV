bind zadaci zadaci_checker c0(.clk(clk), .rst(rst), 
							  .rt_1(rt_1), .rdy_1(rdy_1), .start_1(start_1), .endd_1(endd_1),
							  .er_2(er_2),
							  .er_3(er_3), .rdy_3(rdy_3),
							  .rdy_4(rdy_4), .start_4(start_4),
							  .endd_5(endd_5), .stop_5(stop_5), .er_5(er_5),.rdy_5(rdy_5), .start_5(start_5),
							  .endd_6(endd_6), .stop_6(stop_6), .er_6(er_6), .rdy_6(rdy_6),
							  .endd_7(endd_7), .start_7(start_7), .status_valid_7(status_valid_7), .instartsv_7(instartsv_7),
							  .rt_8(rt_8), .enable_8(enable_8),
							  .rdy_9(rdy_9), .start_9(start_9), .interrupt_9(interrupt_9),
							  .ack_10(ack_10), .req_10(req_10)
							 );
							  
